-- Copyright (C) 1991-2012 Altera Corporation
-- Your use of Altera Corporation's design tools, logic functions 
-- and other software and tools, and its AMPP partner logic 
-- functions, and any output files from any of the foregoing 
-- (including device programming or simulation files), and any 
-- associated documentation or information are expressly subject 
-- to the terms and conditions of the Altera Program License 
-- Subscription Agreement, Altera MegaCore Function License 
-- Agreement, or other applicable license agreement, including, 
-- without limitation, that your use is for the sole purpose of 
-- programming logic devices manufactured by Altera and sold by 
-- Altera or its authorized distributors.  Please refer to the 
-- applicable agreement for further details.

-- PROGRAM		"Quartus II 32-bit"
-- VERSION		"Version 12.1 Build 177 11/07/2012 SJ Full Version"
-- CREATED		"Mon Oct 30 22:14:29 2017"

LIBRARY ieee;
USE ieee.std_logic_1164.all; 

LIBRARY work;

ENTITY display IS 
	PORT
	(
		A :  IN  STD_LOGIC;
		B :  IN  STD_LOGIC;
		C :  IN  STD_LOGIC;
		D :  IN  STD_LOGIC;
		LU :  OUT  STD_LOGIC;
		RU :  OUT  STD_LOGIC;
		RL :  OUT  STD_LOGIC;
		MU :  OUT  STD_LOGIC;
		MM :  OUT  STD_LOGIC;
		ML :  OUT  STD_LOGIC;
		LL :  OUT  STD_LOGIC
	);
END display;

ARCHITECTURE bdf_type OF display IS 

SIGNAL	NA :  STD_LOGIC;
SIGNAL	NB :  STD_LOGIC;
SIGNAL	NC :  STD_LOGIC;
SIGNAL	ND :  STD_LOGIC;
SIGNAL	NLL :  STD_LOGIC;
SIGNAL	NLU :  STD_LOGIC;
SIGNAL	NML :  STD_LOGIC;
SIGNAL	NMM :  STD_LOGIC;
SIGNAL	NMU :  STD_LOGIC;
SIGNAL	NRL :  STD_LOGIC;
SIGNAL	NRU :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_0 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_1 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_2 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_3 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_4 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_5 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_6 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_7 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_8 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_9 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_10 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_11 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_12 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_13 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_14 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_15 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_16 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_17 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_18 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_19 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_20 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_21 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_22 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_23 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_24 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_25 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_26 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_27 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_28 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_29 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_30 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_31 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_32 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_33 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_34 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_35 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_36 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_37 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_38 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_39 :  STD_LOGIC;


BEGIN 
SYNTHESIZED_WIRE_5 <= '0';
SYNTHESIZED_WIRE_15 <= '0';
SYNTHESIZED_WIRE_23 <= '0';
SYNTHESIZED_WIRE_29 <= '0';
SYNTHESIZED_WIRE_35 <= '0';






NA <= NOT(A);



SYNTHESIZED_WIRE_0 <= NB AND C;


SYNTHESIZED_WIRE_2 <= C AND ND;


SYNTHESIZED_WIRE_1 <= A AND NB;


SYNTHESIZED_WIRE_3 <= A AND D;


SYNTHESIZED_WIRE_6 <= NB AND ND;


SYNTHESIZED_WIRE_8 <= NA AND C;


SYNTHESIZED_WIRE_7 <= B AND C;


NB <= NOT(B);



SYNTHESIZED_WIRE_9 <= A AND ND;


SYNTHESIZED_WIRE_12 <= NA AND NB;


SYNTHESIZED_WIRE_14 <= NB AND ND;


SYNTHESIZED_WIRE_18 <= NA AND NC;


SYNTHESIZED_WIRE_20 <= NA AND D;


SYNTHESIZED_WIRE_19 <= NC AND D;


SYNTHESIZED_WIRE_21 <= NA AND B;


SYNTHESIZED_WIRE_22 <= A AND NB;


NC <= NOT(C);



SYNTHESIZED_WIRE_25 <= A AND NB;


SYNTHESIZED_WIRE_4 <= NA AND B AND NC;


SYNTHESIZED_WIRE_10 <= NA AND B AND D;


SYNTHESIZED_WIRE_11 <= A AND NB AND NC;


SYNTHESIZED_WIRE_17 <= NA AND C AND D;


SYNTHESIZED_WIRE_24 <= NC AND ND;


SYNTHESIZED_WIRE_26 <= B AND ND;


SYNTHESIZED_WIRE_27 <= A AND C;


ND <= NOT(D);



SYNTHESIZED_WIRE_28 <= NA AND B AND NC;


SYNTHESIZED_WIRE_36 <= NB AND ND;


SYNTHESIZED_WIRE_39 <= C AND ND;


SYNTHESIZED_WIRE_37 <= A AND C;


SYNTHESIZED_WIRE_38 <= A AND B;


SYNTHESIZED_WIRE_30 <= NA AND NB AND ND;


SYNTHESIZED_WIRE_32 <= NB AND C AND D;


SYNTHESIZED_WIRE_31 <= B AND NC AND D;


SYNTHESIZED_WIRE_33 <= B AND C AND ND;


SYNTHESIZED_WIRE_34 <= A AND NC AND ND;


NMM <= SYNTHESIZED_WIRE_0 OR SYNTHESIZED_WIRE_1 OR SYNTHESIZED_WIRE_2 OR SYNTHESIZED_WIRE_3 OR SYNTHESIZED_WIRE_4 OR SYNTHESIZED_WIRE_5;


NMU <= SYNTHESIZED_WIRE_6 OR SYNTHESIZED_WIRE_7 OR SYNTHESIZED_WIRE_8 OR SYNTHESIZED_WIRE_9 OR SYNTHESIZED_WIRE_10 OR SYNTHESIZED_WIRE_11;


NRU <= SYNTHESIZED_WIRE_12 OR SYNTHESIZED_WIRE_13 OR SYNTHESIZED_WIRE_14 OR SYNTHESIZED_WIRE_15 OR SYNTHESIZED_WIRE_16 OR SYNTHESIZED_WIRE_17;


NRL <= SYNTHESIZED_WIRE_18 OR SYNTHESIZED_WIRE_19 OR SYNTHESIZED_WIRE_20 OR SYNTHESIZED_WIRE_21 OR SYNTHESIZED_WIRE_22 OR SYNTHESIZED_WIRE_23;


NLU <= SYNTHESIZED_WIRE_24 OR SYNTHESIZED_WIRE_25 OR SYNTHESIZED_WIRE_26 OR SYNTHESIZED_WIRE_27 OR SYNTHESIZED_WIRE_28 OR SYNTHESIZED_WIRE_29;


NML <= SYNTHESIZED_WIRE_30 OR SYNTHESIZED_WIRE_31 OR SYNTHESIZED_WIRE_32 OR SYNTHESIZED_WIRE_33 OR SYNTHESIZED_WIRE_34 OR SYNTHESIZED_WIRE_35;


NLL <= SYNTHESIZED_WIRE_36 OR SYNTHESIZED_WIRE_37 OR SYNTHESIZED_WIRE_38 OR SYNTHESIZED_WIRE_39;


LU <= NOT(NLU);



RU <= NOT(NRU);



RL <= NOT(NRL);



MU <= NOT(NMU);



MM <= NOT(NMM);



ML <= NOT(NML);



SYNTHESIZED_WIRE_16 <= NC AND NA AND ND;




SYNTHESIZED_WIRE_13 <= A AND D AND NC;


LL <= NOT(NLL);



END bdf_type;